module parser()
    
endmodule