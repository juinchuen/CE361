// Testbench for Northwestern - CompEng 361 - Lab2
`include "pipelined_cpu.v"

module tb;
    reg clk, rst;
    reg exit;
    wire halt;
    

    // Single Cycle CPU instantiation
    PipelinedCPU CPU (halt, clk,rst);

    // Clock Period = 10 time units
    always
        #5 clk = ~clk;

    always @(posedge clk)
        if (halt)
        exit = 1;
   
    initial begin
        $dumpfile("pipelined_cpu.vcd");
        $dumpvars(0, tb);
        $display("Test Bench for pipelined_cpu\n");
        // Clock and reset steup
        #0 rst = 1; clk = 0; exit =0;
        #0 rst = 0;
        #0 rst = 1;

        // Load program
        #0 $readmemh("mem_in.hex", CPU.IMEM.Mem);
        #0 $readmemh("mem_in.hex", CPU.DMEM.Mem);
        #0 $readmemh("regs_in.hex", CPU.RF.Mem);

        // Feel free to modify to inspect whatever you want
        #0 $monitor($time,, "PC=%08x IR=%08x halt=%x exit=%x", CPU.PC, CPU.InstWord, halt, exit);

        // Exit???
        wait(exit);
        
        // Dump registers
        #0 $writememh("regs_out.hex", CPU.RF.Mem);

        // Dump memory
        #0 $writememh("mem_out.hex", CPU.DMEM.Mem);

        $finish;      
    end
   

endmodule // tb

