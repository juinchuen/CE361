module parser()

endmodule